/**
 * NOTE: you should not need to change this file! This file will be swapped out for a grading
 * "skeleton" for testing. We will also remove your imem and dmem file.
 *
 * NOTE: skeleton should be your top-level module!
 *
 * This skeleton file serves as a wrapper around the processor to provide certain control signals
 * and interfaces to memory elements. This structure allows for easier testing, as it is easier to
 * inspect which signals the processor tries to assert when.
 */

module skeleton(clock, reset,
//for testing
  data_writeReg, ctrl_writeEnable, ctrl_writeReg, wren, address_dmem, data, ctrl_readRegA, 
  ctrl_readRegB, address_imem, flush_overall, opcode, control, control_prev, reg3, signal_to_write
);
    input clock, reset;
	 
    output [11:0] address_imem;
	 output flush_overall;
	 output[31:0] control;
	 output[31:0] control_prev;
    wire [31:0] q_imem;
	 output [4:0] opcode;
	 assign opcode = q_imem[31:27];
    imem my_imem(
        .address    (address_imem),            // address of data
        .clock      (~clock),                  // you may need to invert the clock
        .q          (q_imem)                   // the raw instruction
    );

    /** DMEM **/
    // Figure out how to generate a Quartus syncram component and commit the generated verilog file.
    // Make sure you configure it correctly!
    //wire [11:0] address_dmem;
    //wire [31:0] data;
   // wire wren;
    wire [31:0] q_dmem; //uncomment
	 
	 //DELETE
	 
	 output [31:0] data_writeReg;
	 output ctrl_writeEnable, wren;
	 output [4:0] ctrl_writeReg;
	 
	 output [11:0] address_dmem;
    output [31:0] data;
	 output [4:0]  ctrl_readRegA, ctrl_readRegB;
	 
	 
	 //END DELETE
	 
	 
	 
	 
	 
    dmem my_dmem(
        .address    (address_dmem),       // address of data
        .clock      (~clock),                  // may need to invert the clock
        .data	    (data),    // data you want to write
        .wren	    (wren),      // write enable
        .q          (q_dmem)    // data from dmem
    );

    /** REGFILE **/
    // Instantiate your regfile
	 //uncomment these 
		// wire ctrl_writeEnable;
		//wire [4:0] ctrl_writeReg
		// wire [4:0]  ctrl_readRegA, ctrl_readRegB;
		// wire [31:0] data_writeReg;
    wire [31:0] data_readRegA, data_readRegB;
	 
	 output[31:0] reg3; //for notes 
	 input signal_to_write; //will be sent from the display
    regfile my_regfile(
        clock,
        ctrl_writeEnable,
        reset,
        ctrl_writeReg,
        ctrl_readRegA,
        ctrl_readRegB,
        data_writeReg,
        data_readRegA,
        data_readRegB,
		  reg3,
		  signal_to_write //r1 will be written high if the game needs a new note
    );

    /** PROCESSOR **/
    processor my_processor(
        // Control signals
        clock,                          // I: The master clock
        reset,                          // I: A reset signal

        // Imem
        address_imem,                   // O: The address of the data to get from imem
        q_imem,                         // I: The data from imem
 
        // Dmem
        address_dmem,                   // O: The address of the data to get or put from/to dmem
        data,                           // O: The data to write to dmem
        wren,                           // O: Write enable for dmem
        q_dmem,                         // I: The data from dmem

        // Regfile
        ctrl_writeEnable,               // O: Write enable for regfile
        ctrl_writeReg,                  // O: Register to write to in regfile
        ctrl_readRegA,                  // O: Register to read from port A of regfile
        ctrl_readRegB,                  // O: Register to read from port B of regfile
        data_writeReg,                  // O: Data to write to for regfile
        data_readRegA,                  // I: Data from port A of regfile
        data_readRegB, 						  // I: Data from port B of regfile
		  //read_3,
   flush_overall, control, control_prev
	 );

endmodule
